// Hello World en Verilog

module hello;
  initial
    begin
      $display("Hello, World");
      $display("I am an Icarus Verilog Program.");
      $finish ;
    end
endmodule
